module div(
    input x,
    output divx
);
    assign divx = x / 4'd10;

endmodule // div