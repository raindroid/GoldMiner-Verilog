/**
 *  this module is used to manipulate the ram
 *  and ideally avoid conflict and make life easier
 **/

module MapMan(
    input clock, resetn,
    input 
);
    

endmodule // MapManip