module index(
  
);
    
endmodule // index