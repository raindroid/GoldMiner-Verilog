
//To access data (signX[degree/2] ? -1 : 1) * absX[degree / 2 * 10 + 9 : degree / 2 * 10] / 100
module trigonometry(
    input clock, enable,
    inout [1799: 0] absX, absY,
    inout [179:0] signX, signY
);

integer [1799: 0] rx, ry;
integer [180:0] rsx, rsy;
assign absX = rx;
assign absY = ry;
assign signX = rsx;
assign signY = rsy;

always @(posedge clock) begin
    if (enable) begin //start init our big big table


		rx[1799:1790]	= 10'd 99;
		ry[1799:1790]	= 10'd  3;
		rsx[179]  	= 1'b   0;
		rsy[179]  	= 1'b   1;
		rx[1789:1780]	= 10'd 99;
		ry[1789:1780]	= 10'd  6;
		rsx[178]  	= 1'b   0;
		rsy[178]  	= 1'b   1;
		rx[1779:1770]	= 10'd 99;
		ry[1779:1770]	= 10'd 10;
		rsx[177]  	= 1'b   0;
		rsy[177]  	= 1'b   1;
		rx[1769:1760]	= 10'd 99;
		ry[1769:1760]	= 10'd 13;
		rsx[176]  	= 1'b   0;
		rsy[176]  	= 1'b   1;
		rx[1759:1750]	= 10'd 98;
		ry[1759:1750]	= 10'd 17;
		rsx[175]  	= 1'b   0;
		rsy[175]  	= 1'b   1;
		rx[1749:1740]	= 10'd 97;
		ry[1749:1740]	= 10'd 20;
		rsx[174]  	= 1'b   0;
		rsy[174]  	= 1'b   1;
		rx[1739:1730]	= 10'd 97;
		ry[1739:1730]	= 10'd 24;
		rsx[173]  	= 1'b   0;
		rsy[173]  	= 1'b   1;
		rx[1729:1720]	= 10'd 96;
		ry[1729:1720]	= 10'd 27;
		rsx[172]  	= 1'b   0;
		rsy[172]  	= 1'b   1;
		rx[1719:1710]	= 10'd 95;
		ry[1719:1710]	= 10'd 30;
		rsx[171]  	= 1'b   0;
		rsy[171]  	= 1'b   1;
		rx[1709:1700]	= 10'd 93;
		ry[1709:1700]	= 10'd 34;
		rsx[170]  	= 1'b   0;
		rsy[170]  	= 1'b   1;
		rx[1699:1690]	= 10'd 92;
		ry[1699:1690]	= 10'd 37;
		rsx[169]  	= 1'b   0;
		rsy[169]  	= 1'b   1;
		rx[1689:1680]	= 10'd 91;
		ry[1689:1680]	= 10'd 40;
		rsx[168]  	= 1'b   0;
		rsy[168]  	= 1'b   1;
		rx[1679:1670]	= 10'd 89;
		ry[1679:1670]	= 10'd 43;
		rsx[167]  	= 1'b   0;
		rsy[167]  	= 1'b   1;
		rx[1669:1660]	= 10'd 88;
		ry[1669:1660]	= 10'd 46;
		rsx[166]  	= 1'b   0;
		rsy[166]  	= 1'b   1;
		rx[1659:1650]	= 10'd 86;
		ry[1659:1650]	= 10'd 50;
		rsx[165]  	= 1'b   0;
		rsy[165]  	= 1'b   1;
		rx[1649:1640]	= 10'd 84;
		ry[1649:1640]	= 10'd 52;
		rsx[164]  	= 1'b   0;
		rsy[164]  	= 1'b   1;
		rx[1639:1630]	= 10'd 82;
		ry[1639:1630]	= 10'd 55;
		rsx[163]  	= 1'b   0;
		rsy[163]  	= 1'b   1;
		rx[1629:1620]	= 10'd 80;
		ry[1629:1620]	= 10'd 58;
		rsx[162]  	= 1'b   0;
		rsy[162]  	= 1'b   1;
		rx[1619:1610]	= 10'd 78;
		ry[1619:1610]	= 10'd 61;
		rsx[161]  	= 1'b   0;
		rsy[161]  	= 1'b   1;
		rx[1609:1600]	= 10'd 76;
		ry[1609:1600]	= 10'd 64;
		rsx[160]  	= 1'b   0;
		rsy[160]  	= 1'b   1;
		rx[1599:1590]	= 10'd 74;
		ry[1599:1590]	= 10'd 66;
		rsx[159]  	= 1'b   0;
		rsy[159]  	= 1'b   1;
		rx[1589:1580]	= 10'd 71;
		ry[1589:1580]	= 10'd 69;
		rsx[158]  	= 1'b   0;
		rsy[158]  	= 1'b   1;
		rx[1579:1570]	= 10'd 69;
		ry[1579:1570]	= 10'd 71;
		rsx[157]  	= 1'b   0;
		rsy[157]  	= 1'b   1;
		rx[1569:1560]	= 10'd 66;
		ry[1569:1560]	= 10'd 74;
		rsx[156]  	= 1'b   0;
		rsy[156]  	= 1'b   1;
		rx[1559:1550]	= 10'd 64;
		ry[1559:1550]	= 10'd 76;
		rsx[155]  	= 1'b   0;
		rsy[155]  	= 1'b   1;
		rx[1549:1540]	= 10'd 61;
		ry[1549:1540]	= 10'd 78;
		rsx[154]  	= 1'b   0;
		rsy[154]  	= 1'b   1;
		rx[1539:1530]	= 10'd 58;
		ry[1539:1530]	= 10'd 80;
		rsx[153]  	= 1'b   0;
		rsy[153]  	= 1'b   1;
		rx[1529:1520]	= 10'd 55;
		ry[1529:1520]	= 10'd 82;
		rsx[152]  	= 1'b   0;
		rsy[152]  	= 1'b   1;
		rx[1519:1510]	= 10'd 52;
		ry[1519:1510]	= 10'd 84;
		rsx[151]  	= 1'b   0;
		rsy[151]  	= 1'b   1;
		rx[1509:1500]	= 10'd 50;
		ry[1509:1500]	= 10'd 86;
		rsx[150]  	= 1'b   0;
		rsy[150]  	= 1'b   1;
		rx[1499:1490]	= 10'd 46;
		ry[1499:1490]	= 10'd 88;
		rsx[149]  	= 1'b   0;
		rsy[149]  	= 1'b   1;
		rx[1489:1480]	= 10'd 43;
		ry[1489:1480]	= 10'd 89;
		rsx[148]  	= 1'b   0;
		rsy[148]  	= 1'b   1;
		rx[1479:1470]	= 10'd 40;
		ry[1479:1470]	= 10'd 91;
		rsx[147]  	= 1'b   0;
		rsy[147]  	= 1'b   1;
		rx[1469:1460]	= 10'd 37;
		ry[1469:1460]	= 10'd 92;
		rsx[146]  	= 1'b   0;
		rsy[146]  	= 1'b   1;
		rx[1459:1450]	= 10'd 34;
		ry[1459:1450]	= 10'd 93;
		rsx[145]  	= 1'b   0;
		rsy[145]  	= 1'b   1;
		rx[1449:1440]	= 10'd 30;
		ry[1449:1440]	= 10'd 95;
		rsx[144]  	= 1'b   0;
		rsy[144]  	= 1'b   1;
		rx[1439:1430]	= 10'd 27;
		ry[1439:1430]	= 10'd 96;
		rsx[143]  	= 1'b   0;
		rsy[143]  	= 1'b   1;
		rx[1429:1420]	= 10'd 24;
		ry[1429:1420]	= 10'd 97;
		rsx[142]  	= 1'b   0;
		rsy[142]  	= 1'b   1;
		rx[1419:1410]	= 10'd 20;
		ry[1419:1410]	= 10'd 97;
		rsx[141]  	= 1'b   0;
		rsy[141]  	= 1'b   1;
		rx[1409:1400]	= 10'd 17;
		ry[1409:1400]	= 10'd 98;
		rsx[140]  	= 1'b   0;
		rsy[140]  	= 1'b   1;
		rx[1399:1390]	= 10'd 13;
		ry[1399:1390]	= 10'd 99;
		rsx[139]  	= 1'b   0;
		rsy[139]  	= 1'b   1;
		rx[1389:1380]	= 10'd 10;
		ry[1389:1380]	= 10'd 99;
		rsx[138]  	= 1'b   0;
		rsy[138]  	= 1'b   1;
		rx[1379:1370]	= 10'd  6;
		ry[1379:1370]	= 10'd 99;
		rsx[137]  	= 1'b   0;
		rsy[137]  	= 1'b   1;
		rx[1369:1360]	= 10'd  3;
		ry[1369:1360]	= 10'd 99;
		rsx[136]  	= 1'b   0;
		rsy[136]  	= 1'b   1;
		rx[1359:1350]	= 10'd  0;
		ry[1359:1350]	= 10'd100;
		rsx[135]  	= 1'b   0;
		rsy[135]  	= 1'b   1;
		rx[1349:1340]	= 10'd  3;
		ry[1349:1340]	= 10'd 99;
		rsx[134]  	= 1'b   1;
		rsy[134]  	= 1'b   1;
		rx[1339:1330]	= 10'd  6;
		ry[1339:1330]	= 10'd 99;
		rsx[133]  	= 1'b   1;
		rsy[133]  	= 1'b   1;
		rx[1329:1320]	= 10'd 10;
		ry[1329:1320]	= 10'd 99;
		rsx[132]  	= 1'b   1;
		rsy[132]  	= 1'b   1;
		rx[1319:1310]	= 10'd 13;
		ry[1319:1310]	= 10'd 99;
		rsx[131]  	= 1'b   1;
		rsy[131]  	= 1'b   1;
		rx[1309:1300]	= 10'd 17;
		ry[1309:1300]	= 10'd 98;
		rsx[130]  	= 1'b   1;
		rsy[130]  	= 1'b   1;
		rx[1299:1290]	= 10'd 20;
		ry[1299:1290]	= 10'd 97;
		rsx[129]  	= 1'b   1;
		rsy[129]  	= 1'b   1;
		rx[1289:1280]	= 10'd 24;
		ry[1289:1280]	= 10'd 97;
		rsx[128]  	= 1'b   1;
		rsy[128]  	= 1'b   1;
		rx[1279:1270]	= 10'd 27;
		ry[1279:1270]	= 10'd 96;
		rsx[127]  	= 1'b   1;
		rsy[127]  	= 1'b   1;
		rx[1269:1260]	= 10'd 30;
		ry[1269:1260]	= 10'd 95;
		rsx[126]  	= 1'b   1;
		rsy[126]  	= 1'b   1;
		rx[1259:1250]	= 10'd 34;
		ry[1259:1250]	= 10'd 93;
		rsx[125]  	= 1'b   1;
		rsy[125]  	= 1'b   1;
		rx[1249:1240]	= 10'd 37;
		ry[1249:1240]	= 10'd 92;
		rsx[124]  	= 1'b   1;
		rsy[124]  	= 1'b   1;
		rx[1239:1230]	= 10'd 40;
		ry[1239:1230]	= 10'd 91;
		rsx[123]  	= 1'b   1;
		rsy[123]  	= 1'b   1;
		rx[1229:1220]	= 10'd 43;
		ry[1229:1220]	= 10'd 89;
		rsx[122]  	= 1'b   1;
		rsy[122]  	= 1'b   1;
		rx[1219:1210]	= 10'd 46;
		ry[1219:1210]	= 10'd 88;
		rsx[121]  	= 1'b   1;
		rsy[121]  	= 1'b   1;
		rx[1209:1200]	= 10'd 50;
		ry[1209:1200]	= 10'd 86;
		rsx[120]  	= 1'b   1;
		rsy[120]  	= 1'b   1;
		rx[1199:1190]	= 10'd 52;
		ry[1199:1190]	= 10'd 84;
		rsx[119]  	= 1'b   1;
		rsy[119]  	= 1'b   1;
		rx[1189:1180]	= 10'd 55;
		ry[1189:1180]	= 10'd 82;
		rsx[118]  	= 1'b   1;
		rsy[118]  	= 1'b   1;
		rx[1179:1170]	= 10'd 58;
		ry[1179:1170]	= 10'd 80;
		rsx[117]  	= 1'b   1;
		rsy[117]  	= 1'b   1;
		rx[1169:1160]	= 10'd 61;
		ry[1169:1160]	= 10'd 78;
		rsx[116]  	= 1'b   1;
		rsy[116]  	= 1'b   1;
		rx[1159:1150]	= 10'd 64;
		ry[1159:1150]	= 10'd 76;
		rsx[115]  	= 1'b   1;
		rsy[115]  	= 1'b   1;
		rx[1149:1140]	= 10'd 66;
		ry[1149:1140]	= 10'd 74;
		rsx[114]  	= 1'b   1;
		rsy[114]  	= 1'b   1;
		rx[1139:1130]	= 10'd 69;
		ry[1139:1130]	= 10'd 71;
		rsx[113]  	= 1'b   1;
		rsy[113]  	= 1'b   1;
		rx[1129:1120]	= 10'd 71;
		ry[1129:1120]	= 10'd 69;
		rsx[112]  	= 1'b   1;
		rsy[112]  	= 1'b   1;
		rx[1119:1110]	= 10'd 74;
		ry[1119:1110]	= 10'd 66;
		rsx[111]  	= 1'b   1;
		rsy[111]  	= 1'b   1;
		rx[1109:1100]	= 10'd 76;
		ry[1109:1100]	= 10'd 64;
		rsx[110]  	= 1'b   1;
		rsy[110]  	= 1'b   1;
		rx[1099:1090]	= 10'd 78;
		ry[1099:1090]	= 10'd 61;
		rsx[109]  	= 1'b   1;
		rsy[109]  	= 1'b   1;
		rx[1089:1080]	= 10'd 80;
		ry[1089:1080]	= 10'd 58;
		rsx[108]  	= 1'b   1;
		rsy[108]  	= 1'b   1;
		rx[1079:1070]	= 10'd 82;
		ry[1079:1070]	= 10'd 55;
		rsx[107]  	= 1'b   1;
		rsy[107]  	= 1'b   1;
		rx[1069:1060]	= 10'd 84;
		ry[1069:1060]	= 10'd 52;
		rsx[106]  	= 1'b   1;
		rsy[106]  	= 1'b   1;
		rx[1059:1050]	= 10'd 86;
		ry[1059:1050]	= 10'd 50;
		rsx[105]  	= 1'b   1;
		rsy[105]  	= 1'b   1;
		rx[1049:1040]	= 10'd 88;
		ry[1049:1040]	= 10'd 46;
		rsx[104]  	= 1'b   1;
		rsy[104]  	= 1'b   1;
		rx[1039:1030]	= 10'd 89;
		ry[1039:1030]	= 10'd 43;
		rsx[103]  	= 1'b   1;
		rsy[103]  	= 1'b   1;
		rx[1029:1020]	= 10'd 91;
		ry[1029:1020]	= 10'd 40;
		rsx[102]  	= 1'b   1;
		rsy[102]  	= 1'b   1;
		rx[1019:1010]	= 10'd 92;
		ry[1019:1010]	= 10'd 37;
		rsx[101]  	= 1'b   1;
		rsy[101]  	= 1'b   1;
		rx[1009:1000]	= 10'd 93;
		ry[1009:1000]	= 10'd 34;
		rsx[100]  	= 1'b   1;
		rsy[100]  	= 1'b   1;
		rx[999:990]	= 10'd 95;
		ry[999:990]	= 10'd 30;
		rsx[99]  	= 1'b   1;
		rsy[99]  	= 1'b   1;
		rx[989:980]	= 10'd 96;
		ry[989:980]	= 10'd 27;
		rsx[98]  	= 1'b   1;
		rsy[98]  	= 1'b   1;
		rx[979:970]	= 10'd 97;
		ry[979:970]	= 10'd 24;
		rsx[97]  	= 1'b   1;
		rsy[97]  	= 1'b   1;
		rx[969:960]	= 10'd 97;
		ry[969:960]	= 10'd 20;
		rsx[96]  	= 1'b   1;
		rsy[96]  	= 1'b   1;
		rx[959:950]	= 10'd 98;
		ry[959:950]	= 10'd 17;
		rsx[95]  	= 1'b   1;
		rsy[95]  	= 1'b   1;
		rx[949:940]	= 10'd 99;
		ry[949:940]	= 10'd 13;
		rsx[94]  	= 1'b   1;
		rsy[94]  	= 1'b   1;
		rx[939:930]	= 10'd 99;
		ry[939:930]	= 10'd 10;
		rsx[93]  	= 1'b   1;
		rsy[93]  	= 1'b   1;
		rx[929:920]	= 10'd 99;
		ry[929:920]	= 10'd  6;
		rsx[92]  	= 1'b   1;
		rsy[92]  	= 1'b   1;
		rx[919:910]	= 10'd 99;
		ry[919:910]	= 10'd  3;
		rsx[91]  	= 1'b   1;
		rsy[91]  	= 1'b   1;
		rx[909:900]	= 10'd100;
		ry[909:900]	= 10'd  0;
		rsx[90]  	= 1'b   1;
		rsy[90]  	= 1'b   0;
		rx[899:890]	= 10'd 99;
		ry[899:890]	= 10'd  3;
		rsx[89]  	= 1'b   1;
		rsy[89]  	= 1'b   0;
		rx[889:880]	= 10'd 99;
		ry[889:880]	= 10'd  6;
		rsx[88]  	= 1'b   1;
		rsy[88]  	= 1'b   0;
		rx[879:870]	= 10'd 99;
		ry[879:870]	= 10'd 10;
		rsx[87]  	= 1'b   1;
		rsy[87]  	= 1'b   0;
		rx[869:860]	= 10'd 99;
		ry[869:860]	= 10'd 13;
		rsx[86]  	= 1'b   1;
		rsy[86]  	= 1'b   0;
		rx[859:850]	= 10'd 98;
		ry[859:850]	= 10'd 17;
		rsx[85]  	= 1'b   1;
		rsy[85]  	= 1'b   0;
		rx[849:840]	= 10'd 97;
		ry[849:840]	= 10'd 20;
		rsx[84]  	= 1'b   1;
		rsy[84]  	= 1'b   0;
		rx[839:830]	= 10'd 97;
		ry[839:830]	= 10'd 24;
		rsx[83]  	= 1'b   1;
		rsy[83]  	= 1'b   0;
		rx[829:820]	= 10'd 96;
		ry[829:820]	= 10'd 27;
		rsx[82]  	= 1'b   1;
		rsy[82]  	= 1'b   0;
		rx[819:810]	= 10'd 95;
		ry[819:810]	= 10'd 30;
		rsx[81]  	= 1'b   1;
		rsy[81]  	= 1'b   0;
		rx[809:800]	= 10'd 93;
		ry[809:800]	= 10'd 34;
		rsx[80]  	= 1'b   1;
		rsy[80]  	= 1'b   0;
		rx[799:790]	= 10'd 92;
		ry[799:790]	= 10'd 37;
		rsx[79]  	= 1'b   1;
		rsy[79]  	= 1'b   0;
		rx[789:780]	= 10'd 91;
		ry[789:780]	= 10'd 40;
		rsx[78]  	= 1'b   1;
		rsy[78]  	= 1'b   0;
		rx[779:770]	= 10'd 89;
		ry[779:770]	= 10'd 43;
		rsx[77]  	= 1'b   1;
		rsy[77]  	= 1'b   0;
		rx[769:760]	= 10'd 88;
		ry[769:760]	= 10'd 46;
		rsx[76]  	= 1'b   1;
		rsy[76]  	= 1'b   0;
		rx[759:750]	= 10'd 86;
		ry[759:750]	= 10'd 49;
		rsx[75]  	= 1'b   1;
		rsy[75]  	= 1'b   0;
		rx[749:740]	= 10'd 84;
		ry[749:740]	= 10'd 52;
		rsx[74]  	= 1'b   1;
		rsy[74]  	= 1'b   0;
		rx[739:730]	= 10'd 82;
		ry[739:730]	= 10'd 55;
		rsx[73]  	= 1'b   1;
		rsy[73]  	= 1'b   0;
		rx[729:720]	= 10'd 80;
		ry[729:720]	= 10'd 58;
		rsx[72]  	= 1'b   1;
		rsy[72]  	= 1'b   0;
		rx[719:710]	= 10'd 78;
		ry[719:710]	= 10'd 61;
		rsx[71]  	= 1'b   1;
		rsy[71]  	= 1'b   0;
		rx[709:700]	= 10'd 76;
		ry[709:700]	= 10'd 64;
		rsx[70]  	= 1'b   1;
		rsy[70]  	= 1'b   0;
		rx[699:690]	= 10'd 74;
		ry[699:690]	= 10'd 66;
		rsx[69]  	= 1'b   1;
		rsy[69]  	= 1'b   0;
		rx[689:680]	= 10'd 71;
		ry[689:680]	= 10'd 69;
		rsx[68]  	= 1'b   1;
		rsy[68]  	= 1'b   0;
		rx[679:670]	= 10'd 69;
		ry[679:670]	= 10'd 71;
		rsx[67]  	= 1'b   1;
		rsy[67]  	= 1'b   0;
		rx[669:660]	= 10'd 66;
		ry[669:660]	= 10'd 74;
		rsx[66]  	= 1'b   1;
		rsy[66]  	= 1'b   0;
		rx[659:650]	= 10'd 64;
		ry[659:650]	= 10'd 76;
		rsx[65]  	= 1'b   1;
		rsy[65]  	= 1'b   0;
		rx[649:640]	= 10'd 61;
		ry[649:640]	= 10'd 78;
		rsx[64]  	= 1'b   1;
		rsy[64]  	= 1'b   0;
		rx[639:630]	= 10'd 58;
		ry[639:630]	= 10'd 80;
		rsx[63]  	= 1'b   1;
		rsy[63]  	= 1'b   0;
		rx[629:620]	= 10'd 55;
		ry[629:620]	= 10'd 82;
		rsx[62]  	= 1'b   1;
		rsy[62]  	= 1'b   0;
		rx[619:610]	= 10'd 52;
		ry[619:610]	= 10'd 84;
		rsx[61]  	= 1'b   1;
		rsy[61]  	= 1'b   0;
		rx[609:600]	= 10'd 49;
		ry[609:600]	= 10'd 86;
		rsx[60]  	= 1'b   1;
		rsy[60]  	= 1'b   0;
		rx[599:590]	= 10'd 46;
		ry[599:590]	= 10'd 88;
		rsx[59]  	= 1'b   1;
		rsy[59]  	= 1'b   0;
		rx[589:580]	= 10'd 43;
		ry[589:580]	= 10'd 89;
		rsx[58]  	= 1'b   1;
		rsy[58]  	= 1'b   0;
		rx[579:570]	= 10'd 40;
		ry[579:570]	= 10'd 91;
		rsx[57]  	= 1'b   1;
		rsy[57]  	= 1'b   0;
		rx[569:560]	= 10'd 37;
		ry[569:560]	= 10'd 92;
		rsx[56]  	= 1'b   1;
		rsy[56]  	= 1'b   0;
		rx[559:550]	= 10'd 34;
		ry[559:550]	= 10'd 93;
		rsx[55]  	= 1'b   1;
		rsy[55]  	= 1'b   0;
		rx[549:540]	= 10'd 30;
		ry[549:540]	= 10'd 95;
		rsx[54]  	= 1'b   1;
		rsy[54]  	= 1'b   0;
		rx[539:530]	= 10'd 27;
		ry[539:530]	= 10'd 96;
		rsx[53]  	= 1'b   1;
		rsy[53]  	= 1'b   0;
		rx[529:520]	= 10'd 24;
		ry[529:520]	= 10'd 97;
		rsx[52]  	= 1'b   1;
		rsy[52]  	= 1'b   0;
		rx[519:510]	= 10'd 20;
		ry[519:510]	= 10'd 97;
		rsx[51]  	= 1'b   1;
		rsy[51]  	= 1'b   0;
		rx[509:500]	= 10'd 17;
		ry[509:500]	= 10'd 98;
		rsx[50]  	= 1'b   1;
		rsy[50]  	= 1'b   0;
		rx[499:490]	= 10'd 13;
		ry[499:490]	= 10'd 99;
		rsx[49]  	= 1'b   1;
		rsy[49]  	= 1'b   0;
		rx[489:480]	= 10'd 10;
		ry[489:480]	= 10'd 99;
		rsx[48]  	= 1'b   1;
		rsy[48]  	= 1'b   0;
		rx[479:470]	= 10'd  6;
		ry[479:470]	= 10'd 99;
		rsx[47]  	= 1'b   1;
		rsy[47]  	= 1'b   0;
		rx[469:460]	= 10'd  3;
		ry[469:460]	= 10'd 99;
		rsx[46]  	= 1'b   1;
		rsy[46]  	= 1'b   0;
		rx[459:450]	= 10'd  0;
		ry[459:450]	= 10'd100;
		rsx[45]  	= 1'b   0;
		rsy[45]  	= 1'b   0;
		rx[449:440]	= 10'd  3;
		ry[449:440]	= 10'd 99;
		rsx[44]  	= 1'b   0;
		rsy[44]  	= 1'b   0;
		rx[439:430]	= 10'd  6;
		ry[439:430]	= 10'd 99;
		rsx[43]  	= 1'b   0;
		rsy[43]  	= 1'b   0;
		rx[429:420]	= 10'd 10;
		ry[429:420]	= 10'd 99;
		rsx[42]  	= 1'b   0;
		rsy[42]  	= 1'b   0;
		rx[419:410]	= 10'd 13;
		ry[419:410]	= 10'd 99;
		rsx[41]  	= 1'b   0;
		rsy[41]  	= 1'b   0;
		rx[409:400]	= 10'd 17;
		ry[409:400]	= 10'd 98;
		rsx[40]  	= 1'b   0;
		rsy[40]  	= 1'b   0;
		rx[399:390]	= 10'd 20;
		ry[399:390]	= 10'd 97;
		rsx[39]  	= 1'b   0;
		rsy[39]  	= 1'b   0;
		rx[389:380]	= 10'd 24;
		ry[389:380]	= 10'd 97;
		rsx[38]  	= 1'b   0;
		rsy[38]  	= 1'b   0;
		rx[379:370]	= 10'd 27;
		ry[379:370]	= 10'd 96;
		rsx[37]  	= 1'b   0;
		rsy[37]  	= 1'b   0;
		rx[369:360]	= 10'd 30;
		ry[369:360]	= 10'd 95;
		rsx[36]  	= 1'b   0;
		rsy[36]  	= 1'b   0;
		rx[359:350]	= 10'd 34;
		ry[359:350]	= 10'd 93;
		rsx[35]  	= 1'b   0;
		rsy[35]  	= 1'b   0;
		rx[349:340]	= 10'd 37;
		ry[349:340]	= 10'd 92;
		rsx[34]  	= 1'b   0;
		rsy[34]  	= 1'b   0;
		rx[339:330]	= 10'd 40;
		ry[339:330]	= 10'd 91;
		rsx[33]  	= 1'b   0;
		rsy[33]  	= 1'b   0;
		rx[329:320]	= 10'd 43;
		ry[329:320]	= 10'd 89;
		rsx[32]  	= 1'b   0;
		rsy[32]  	= 1'b   0;
		rx[319:310]	= 10'd 46;
		ry[319:310]	= 10'd 88;
		rsx[31]  	= 1'b   0;
		rsy[31]  	= 1'b   0;
		rx[309:300]	= 10'd 50;
		ry[309:300]	= 10'd 86;
		rsx[30]  	= 1'b   0;
		rsy[30]  	= 1'b   0;
		rx[299:290]	= 10'd 52;
		ry[299:290]	= 10'd 84;
		rsx[29]  	= 1'b   0;
		rsy[29]  	= 1'b   0;
		rx[289:280]	= 10'd 55;
		ry[289:280]	= 10'd 82;
		rsx[28]  	= 1'b   0;
		rsy[28]  	= 1'b   0;
		rx[279:270]	= 10'd 58;
		ry[279:270]	= 10'd 80;
		rsx[27]  	= 1'b   0;
		rsy[27]  	= 1'b   0;
		rx[269:260]	= 10'd 61;
		ry[269:260]	= 10'd 78;
		rsx[26]  	= 1'b   0;
		rsy[26]  	= 1'b   0;
		rx[259:250]	= 10'd 64;
		ry[259:250]	= 10'd 76;
		rsx[25]  	= 1'b   0;
		rsy[25]  	= 1'b   0;
		rx[249:240]	= 10'd 66;
		ry[249:240]	= 10'd 74;
		rsx[24]  	= 1'b   0;
		rsy[24]  	= 1'b   0;
		rx[239:230]	= 10'd 69;
		ry[239:230]	= 10'd 71;
		rsx[23]  	= 1'b   0;
		rsy[23]  	= 1'b   0;
		rx[229:220]	= 10'd 71;
		ry[229:220]	= 10'd 69;
		rsx[22]  	= 1'b   0;
		rsy[22]  	= 1'b   0;
		rx[219:210]	= 10'd 74;
		ry[219:210]	= 10'd 66;
		rsx[21]  	= 1'b   0;
		rsy[21]  	= 1'b   0;
		rx[209:200]	= 10'd 76;
		ry[209:200]	= 10'd 64;
		rsx[20]  	= 1'b   0;
		rsy[20]  	= 1'b   0;
		rx[199:190]	= 10'd 78;
		ry[199:190]	= 10'd 61;
		rsx[19]  	= 1'b   0;
		rsy[19]  	= 1'b   0;
		rx[189:180]	= 10'd 80;
		ry[189:180]	= 10'd 58;
		rsx[18]  	= 1'b   0;
		rsy[18]  	= 1'b   0;
		rx[179:170]	= 10'd 82;
		ry[179:170]	= 10'd 55;
		rsx[17]  	= 1'b   0;
		rsy[17]  	= 1'b   0;
		rx[169:160]	= 10'd 84;
		ry[169:160]	= 10'd 52;
		rsx[16]  	= 1'b   0;
		rsy[16]  	= 1'b   0;
		rx[159:150]	= 10'd 86;
		ry[159:150]	= 10'd 49;
		rsx[15]  	= 1'b   0;
		rsy[15]  	= 1'b   0;
		rx[149:140]	= 10'd 88;
		ry[149:140]	= 10'd 46;
		rsx[14]  	= 1'b   0;
		rsy[14]  	= 1'b   0;
		rx[139:130]	= 10'd 89;
		ry[139:130]	= 10'd 43;
		rsx[13]  	= 1'b   0;
		rsy[13]  	= 1'b   0;
		rx[129:120]	= 10'd 91;
		ry[129:120]	= 10'd 40;
		rsx[12]  	= 1'b   0;
		rsy[12]  	= 1'b   0;
		rx[119:110]	= 10'd 92;
		ry[119:110]	= 10'd 37;
		rsx[11]  	= 1'b   0;
		rsy[11]  	= 1'b   0;
		rx[109:100]	= 10'd 93;
		ry[109:100]	= 10'd 34;
		rsx[10]  	= 1'b   0;
		rsy[10]  	= 1'b   0;
		rx[99:90]	= 10'd 95;
		ry[99:90]	= 10'd 30;
		rsx[9]  	= 1'b   0;
		rsy[9]  	= 1'b   0;
		rx[89:80]	= 10'd 96;
		ry[89:80]	= 10'd 27;
		rsx[8]  	= 1'b   0;
		rsy[8]  	= 1'b   0;
		rx[79:70]	= 10'd 97;
		ry[79:70]	= 10'd 24;
		rsx[7]  	= 1'b   0;
		rsy[7]  	= 1'b   0;
		rx[69:60]	= 10'd 97;
		ry[69:60]	= 10'd 20;
		rsx[6]  	= 1'b   0;
		rsy[6]  	= 1'b   0;
		rx[59:50]	= 10'd 98;
		ry[59:50]	= 10'd 17;
		rsx[5]  	= 1'b   0;
		rsy[5]  	= 1'b   0;
		rx[49:40]	= 10'd 99;
		ry[49:40]	= 10'd 13;
		rsx[4]  	= 1'b   0;
		rsy[4]  	= 1'b   0;
		rx[39:30]	= 10'd 99;
		ry[39:30]	= 10'd 10;
		rsx[3]  	= 1'b   0;
		rsy[3]  	= 1'b   0;
		rx[29:20]	= 10'd 99;
		ry[29:20]	= 10'd  6;
		rsx[2]  	= 1'b   0;
		rsy[2]  	= 1'b   0;
		rx[19:10]	= 10'd 99;
		ry[19:10]	= 10'd  3;
		rsx[1]  	= 1'b   0;
		rsy[1]  	= 1'b   0;
		rx[9:0] 	= 10'd100;
		ry[9:0] 	= 10'd  0;
		rsx[0]  	= 1'b   0;
		rsy[0]  	= 1'b   0;

    end
end
endmodule